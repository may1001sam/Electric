*** SPICE deck for cell XOR_sim{lay} from library XOR
*** Created on Sun Nov 10, 2024 12:25:45
*** Last revised on Thu Jan 02, 2025 22:36:44
*** Written on Thu Jan 02, 2025 22:38:32 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT XOR__XOR FROM CELL XOR:XOR{lay}
.SUBCKT XOR__XOR A B gnd out vdd
Mnmos@0 net@3 A out gnd N L=0.044U W=0.22U AS=0.036P AD=0.025P PS=0.534U PD=0.561U
Mnmos@1 out net@202 net@3 gnd N L=0.044U W=0.22U AS=0.025P AD=0.036P PS=0.561U PD=0.534U
Mnmos@4 net@3 net@191 gnd gnd N L=0.044U W=0.22U AS=0.14P AD=0.025P PS=1.711U PD=0.561U
Mnmos@5 gnd B net@3 gnd N L=0.044U W=0.22U AS=0.025P AD=0.14P PS=0.561U PD=1.711U
Mnmos@7 gnd A net@191 gnd N L=0.044U W=0.22U AS=0.045P AD=0.14P PS=0.935U PD=1.711U
Mnmos@9 net@202 B gnd gnd N L=0.044U W=0.22U AS=0.14P AD=0.044P PS=1.711U PD=0.924U
Mpmos@0 vdd A net@236 vdd P L=0.044U W=0.44U AS=0.024P AD=0.182P PS=0.55U PD=2.338U
Mpmos@1 net@236 net@202 out vdd P L=0.044U W=0.44U AS=0.036P AD=0.024P PS=0.534U PD=0.55U
Mpmos@4 out net@191 net@240 vdd P L=0.044U W=0.44U AS=0.029P AD=0.036P PS=0.572U PD=0.534U
Mpmos@5 net@240 B vdd vdd P L=0.044U W=0.44U AS=0.182P AD=0.029P PS=2.338U PD=0.572U
Mpmos@6 vdd A net@191 vdd P L=0.044U W=0.44U AS=0.045P AD=0.182P PS=0.935U PD=2.338U
Mpmos@7 net@202 B vdd vdd P L=0.044U W=0.44U AS=0.182P AD=0.044P PS=2.338U PD=0.924U
.ENDS XOR__XOR

*** TOP LEVEL CELL: XOR:XOR_sim{lay}
XXOR@0 A B gnd out vdd XOR__XOR

* Spice Code nodes in cell cell 'XOR:XOR_sim{lay}'
vdd vdd 0 DC 0.95
va A 0 DC pwl 10n 0 20n 0.95 50n 0.95 60n 0 90n 0 100n 0.95 130n 0.95 140n 0 170n 0 180n 0.95
vb B 0 DC pwl 10n 0 20n 0.95 100n 0.95 110n 0
.tran 200n
.include C:\Electric\22nm.txt
.END
