*** SPICE deck for cell 2bit_FA_right_sim{lay} from library 2bit_FA
*** Created on Mon Jan 13, 2025 21:37:24
*** Last revised on Mon Jan 13, 2025 21:42:47
*** Written on Mon Jan 13, 2025 21:42:50 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT _2bit_FA__2bit_FA FROM CELL 2bit_FA:2bit_FA{lay}
.SUBCKT _2bit_FA__2bit_FA A0 A1 B0 B1 c-1 c0 G0 G1 gnd P0 P1 s0 s1 vdd
Mnmos@0 gnd b0 net@3 gnd N L=0.044U W=0.22U AS=0.015P AD=0.161P PS=0.352U PD=1.875U
Mnmos@1 net@3 a0 G0 gnd N L=0.044U W=0.22U AS=0.045P AD=0.015P PS=0.689U PD=0.352U
Mnmos@2 net@14 a0 P0 gnd N L=0.044U W=0.44U AS=0.067P AD=0.047P PS=0.858U PD=0.875U
Mnmos@3 P0 net@22 net@14 gnd N L=0.044U W=0.44U AS=0.047P AD=0.067P PS=0.875U PD=0.858U
Mnmos@4 net@14 net@15 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.047P PS=1.875U PD=0.875U
Mnmos@5 gnd b0 net@14 gnd N L=0.044U W=0.44U AS=0.047P AD=0.161P PS=0.875U PD=1.875U
Mnmos@6 gnd a0 net@15 gnd N L=0.044U W=0.44U AS=0.087P AD=0.161P PS=1.584U PD=1.875U
Mnmos@7 net@22 b0 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.087P PS=1.875U PD=1.584U
Mnmos@8 net@64 P0 s0 gnd N L=0.044U W=0.44U AS=0.067P AD=0.047P PS=0.858U PD=0.875U
Mnmos@9 s0 net@71 net@64 gnd N L=0.044U W=0.44U AS=0.047P AD=0.067P PS=0.875U PD=0.858U
Mnmos@10 net@64 net@65 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.047P PS=1.875U PD=0.875U
Mnmos@11 gnd c-1 net@64 gnd N L=0.044U W=0.44U AS=0.047P AD=0.161P PS=0.875U PD=1.875U
Mnmos@12 gnd P0 net@65 gnd N L=0.044U W=0.44U AS=0.087P AD=0.161P PS=1.584U PD=1.875U
Mnmos@13 net@71 c-1 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.087P PS=1.875U PD=1.584U
Mnmos@14 gnd b1 net@195 gnd N L=0.044U W=0.22U AS=0.015P AD=0.161P PS=0.352U PD=1.875U
Mnmos@15 net@195 a1 G1 gnd N L=0.044U W=0.22U AS=0.045P AD=0.015P PS=0.689U PD=0.352U
Mnmos@16 net@206 a1 P1 gnd N L=0.044U W=0.44U AS=0.067P AD=0.047P PS=0.858U PD=0.875U
Mnmos@17 P1 net@214 net@206 gnd N L=0.044U W=0.44U AS=0.047P AD=0.067P PS=0.875U PD=0.858U
Mnmos@18 net@206 net@207 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.047P PS=1.875U PD=0.875U
Mnmos@19 gnd b1 net@206 gnd N L=0.044U W=0.44U AS=0.047P AD=0.161P PS=0.875U PD=1.875U
Mnmos@20 gnd a1 net@207 gnd N L=0.044U W=0.44U AS=0.087P AD=0.161P PS=1.584U PD=1.875U
Mnmos@21 net@214 b1 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.087P PS=1.875U PD=1.584U
Mnmos@22 net@256 P1 s1 gnd N L=0.044U W=0.44U AS=0.067P AD=0.047P PS=0.858U PD=0.875U
Mnmos@23 s1 net@263 net@256 gnd N L=0.044U W=0.44U AS=0.047P AD=0.067P PS=0.875U PD=0.858U
Mnmos@24 net@256 net@257 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.047P PS=1.875U PD=0.875U
Mnmos@25 gnd c0 net@256 gnd N L=0.044U W=0.44U AS=0.047P AD=0.161P PS=0.875U PD=1.875U
Mnmos@26 gnd P1 net@257 gnd N L=0.044U W=0.44U AS=0.087P AD=0.161P PS=1.584U PD=1.875U
Mnmos@27 net@263 c0 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.087P PS=1.875U PD=1.584U
Mpmos@0 vdd b0 G0 vdd P L=0.044U W=0.44U AS=0.045P AD=0.213P PS=0.689U PD=2.695U
Mpmos@1 G0 a0 vdd vdd P L=0.044U W=0.44U AS=0.213P AD=0.045P PS=2.695U PD=0.689U
Mpmos@2 vdd a0 net@48 vdd P L=0.044U W=0.88U AS=0.053P AD=0.213P PS=1.001U PD=2.695U
Mpmos@3 net@48 net@22 P0 vdd P L=0.044U W=0.88U AS=0.067P AD=0.053P PS=0.858U PD=1.001U
Mpmos@4 P0 net@15 net@51 vdd P L=0.044U W=0.88U AS=0.053P AD=0.067P PS=1.001U PD=0.858U
Mpmos@5 net@51 b0 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.053P PS=2.695U PD=1.001U
Mpmos@6 vdd a0 net@15 vdd P L=0.044U W=0.88U AS=0.087P AD=0.213P PS=1.584U PD=2.695U
Mpmos@7 net@22 b0 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.087P PS=2.695U PD=1.584U
Mpmos@8 vdd P0 net@97 vdd P L=0.044U W=0.88U AS=0.053P AD=0.213P PS=1.001U PD=2.695U
Mpmos@9 net@97 net@71 s0 vdd P L=0.044U W=0.88U AS=0.067P AD=0.053P PS=0.858U PD=1.001U
Mpmos@10 s0 net@65 net@100 vdd P L=0.044U W=0.88U AS=0.053P AD=0.067P PS=1.001U PD=0.858U
Mpmos@11 net@100 c-1 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.053P PS=2.695U PD=1.001U
Mpmos@12 vdd P0 net@65 vdd P L=0.044U W=0.88U AS=0.087P AD=0.213P PS=1.584U PD=2.695U
Mpmos@13 net@71 c-1 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.087P PS=2.695U PD=1.584U
Mpmos@14 vdd b1 G1 vdd P L=0.044U W=0.44U AS=0.045P AD=0.213P PS=0.689U PD=2.695U
Mpmos@15 G1 a1 vdd vdd P L=0.044U W=0.44U AS=0.213P AD=0.045P PS=2.695U PD=0.689U
Mpmos@16 vdd a1 net@240 vdd P L=0.044U W=0.88U AS=0.053P AD=0.213P PS=1.001U PD=2.695U
Mpmos@17 net@240 net@214 P1 vdd P L=0.044U W=0.88U AS=0.067P AD=0.053P PS=0.858U PD=1.001U
Mpmos@18 P1 net@207 net@243 vdd P L=0.044U W=0.88U AS=0.053P AD=0.067P PS=1.001U PD=0.858U
Mpmos@19 net@243 b1 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.053P PS=2.695U PD=1.001U
Mpmos@20 vdd a1 net@207 vdd P L=0.044U W=0.88U AS=0.087P AD=0.213P PS=1.584U PD=2.695U
Mpmos@21 net@214 b1 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.087P PS=2.695U PD=1.584U
Mpmos@22 vdd P1 net@289 vdd P L=0.044U W=0.88U AS=0.053P AD=0.213P PS=1.001U PD=2.695U
Mpmos@23 net@289 net@263 s1 vdd P L=0.044U W=0.88U AS=0.067P AD=0.053P PS=0.858U PD=1.001U
Mpmos@24 s1 net@257 net@292 vdd P L=0.044U W=0.88U AS=0.053P AD=0.067P PS=1.001U PD=0.858U
Mpmos@25 net@292 c0 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.053P PS=2.695U PD=1.001U
Mpmos@26 vdd P1 net@257 vdd P L=0.044U W=0.88U AS=0.087P AD=0.213P PS=1.584U PD=2.695U
Mpmos@27 net@263 c0 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.087P PS=2.695U PD=1.584U
.ENDS _2bit_FA__2bit_FA

*** TOP LEVEL CELL: 2bit_FA:2bit_FA_right_sim{lay}
X_2bit_FA@0 A0 A1 B0 B1 c-1 c0 G0 G1 gnd Po P1 s0 s1 vdd _2bit_FA__2bit_FA

* Spice Code nodes in cell cell '2bit_FA:2bit_FA_right_sim{lay}'
vdd vdd 0 DC 0.95
* 2-bit input A
va0 A0 0 PWL(0n 0 10n 0 12n 0.95 51n 0.95 53n 0 95n 0 97n 0.95 140n 0.95 142n 0 183n 0 185n 0.95)
va1 A1 0 PWL(0n 0.95 10n 0.95 12n 0 51n 0 53n 0.95 95n 0.95 97n 0 140n 0 142n 0.95 183n 0.95 185n 0)
* 2-bit input B
vb0 B0 0 PWL(0n 0 95n 0 97n 0.95)
vb1 B1 0 PWL(0n 0.95 95n 0.95 97n 0)
vc-1 C-1 0 DC 0
vc0 C0 0 DC 0
* Transient analysis
.tran 0 200n
* Include model file
.include C:\Electric\22nm.txt
.END
