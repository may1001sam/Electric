*** SPICE deck for cell 2bit_FA{sch} from library 2bit_FA
*** Created on Mon Jan 13, 2025 18:34:07
*** Last revised on Mon Jan 13, 2025 18:44:32
*** Written on Mon Jan 13, 2025 18:44:39 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT inverter__inv FROM CELL inverter:inv{sch}
.SUBCKT inverter__inv in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.044U W=0.22U
Mpmos@0 vdd in out vdd P L=0.044U W=0.44U
.ENDS inverter__inv

*** SUBCIRCUIT XOR__XOR FROM CELL XOR:XOR{sch}
.SUBCKT XOR__XOR A B out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@8 out A net@13 gnd N L=0.044U W=0.44U
Mnmos@9 out net@57 net@13 gnd N L=0.044U W=0.44U
Mnmos@10 net@13 B gnd gnd N L=0.044U W=0.44U
Mnmos@11 net@13 net@56 gnd gnd N L=0.044U W=0.44U
Mpmos@8 vdd A net@1 vdd P L=0.044U W=0.88U
Mpmos@9 net@1 net@57 out vdd P L=0.044U W=0.88U
Mpmos@10 vdd B net@2 vdd P L=0.044U W=0.88U
Mpmos@11 net@2 net@56 out vdd P L=0.044U W=0.88U
Xinv@0 A net@56 inverter__inv
Xinv@1 B net@57 inverter__inv
.ENDS XOR__XOR

*** SUBCIRCUIT NAND__nand FROM CELL NAND:nand{sch}
.SUBCKT NAND__nand A B out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out A net@11 gnd N L=0.044U W=0.22U
Mnmos@1 net@11 B gnd gnd N L=0.044U W=0.22U
Mpmos@1 vdd A out vdd P L=0.044U W=0.44U
Mpmos@2 vdd B out vdd P L=0.044U W=0.44U
.ENDS NAND__nand

*** SUBCIRCUIT FA_new__FA_new FROM CELL FA_new:FA_new{sch}
.SUBCKT FA_new__FA_new A B Cin G P Sum
** GLOBAL gnd
** GLOBAL vdd
XXOR@0 A B P XOR__XOR
XXOR@1 P Cin Sum XOR__XOR
Xnand@0 A B G NAND__nand
.ENDS FA_new__FA_new

.global gnd vdd

*** TOP LEVEL CELL: 2bit_FA{sch}
XFA_new@0 A1 B1 C0 G1 P1 S1 FA_new__FA_new
XFA_new@1 A0 B0 C-1 G0 P0 S0 FA_new__FA_new

* Spice Code nodes in cell cell '2bit_FA{sch}'
vdd vdd 0 DC 0.95
* 2-bit input A
va0 A0 0 PWL(0n 0 10n 0 12n 0.95 51n 0.95 53n 0 95n 0 97n 0.95 140n 0.95 142n 0 183n 0 185n 0.95)
va1 A1 0 PWL(0n 0.95 10n 0.95 12n 0 51n 0 53n 0.95 95n 0.95 97n 0 140n 0 142n 0.95 183n 0.95 185n 0)
* 2-bit input B
vb0 B0 0 PWL(0n 0 95n 0 97n 0.95)
vb1 B1 0 PWL(0n 0.95 95n 0.95 97n 0)
vc-1 C-1 0 DC 0
vc0 C0 0 DC 0
* Transient analysis
.tran 0 200n
* Include model file
.include C:\Electric\22nm.txt
.END
