*** SPICE deck for cell XOR_sim{lay} from library XOR
*** Created on Sun Nov 10, 2024 12:25:45
*** Last revised on Fri Jan 10, 2025 13:17:34
*** Written on Fri Jan 10, 2025 13:18:09 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT XOR__XOR FROM CELL XOR:XOR{lay}
.SUBCKT XOR__XOR A B gnd out vdd
Mnmos@0 net@3 A out gnd N L=0.044U W=0.44U AS=0.067P AD=0.047P PS=0.858U PD=0.875U
Mnmos@1 out net@256 net@3 gnd N L=0.044U W=0.44U AS=0.047P AD=0.067P PS=0.875U PD=0.858U
Mnmos@4 net@3 net@199 gnd gnd N L=0.044U W=0.44U AS=0.165P AD=0.047P PS=2.04U PD=0.875U
Mnmos@5 gnd B net@3 gnd N L=0.044U W=0.44U AS=0.047P AD=0.165P PS=0.875U PD=2.04U
Mnmos@7 gnd A net@199 gnd N L=0.044U W=0.44U AS=0.087P AD=0.165P PS=1.584U PD=2.04U
Mnmos@9 net@256 B gnd gnd N L=0.044U W=0.44U AS=0.165P AD=0.087P PS=2.04U PD=1.584U
Mpmos@0 vdd A net@477 vdd P L=0.044U W=0.88U AS=0.053P AD=0.238P PS=1.001U PD=3.196U
Mpmos@1 net@477 net@256 out vdd P L=0.044U W=0.88U AS=0.067P AD=0.053P PS=0.858U PD=1.001U
Mpmos@4 out net@199 net@497 vdd P L=0.044U W=0.88U AS=0.053P AD=0.067P PS=1.001U PD=0.858U
Mpmos@5 net@497 B vdd vdd P L=0.044U W=0.88U AS=0.238P AD=0.053P PS=3.196U PD=1.001U
Mpmos@6 vdd A net@199 vdd P L=0.044U W=0.88U AS=0.087P AD=0.238P PS=1.584U PD=3.196U
Mpmos@7 net@256 B vdd vdd P L=0.044U W=0.88U AS=0.238P AD=0.087P PS=3.196U PD=1.584U
.ENDS XOR__XOR

*** TOP LEVEL CELL: XOR:XOR_sim{lay}
XXOR@0 A B gnd out vdd XOR__XOR

* Spice Code nodes in cell cell 'XOR:XOR_sim{lay}'
vdd vdd 0 DC 0.95
va A 0 DC pwl 10n 0 20n 0.95 50n 0.95 60n 0 90n 0 100n 0.95 130n 0.95 140n 0 170n 0 180n 0.95
vb B 0 DC pwl 10n 0 20n 0.95 115n 0.95 120n 0
.tran 200n
.include C:\Electric\22nm.txt
.END
