*** SPICE deck for cell Repeater_sim{lay} from library Repeater
*** Created on Sat Jan 04, 2025 21:13:35
*** Last revised on Sat Jan 04, 2025 21:14:53
*** Written on Sat Jan 04, 2025 21:15:04 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT inverter__inv FROM CELL inverter:inv{lay}
.SUBCKT inverter__inv gnd in out vdd
Mnmos@0 gnd in out gnd N L=0.044U W=0.22U AS=0.058P AD=0.099P PS=1.012U PD=2.112U
Mpmos@0 vdd in out vdd P L=0.044U W=0.44U AS=0.058P AD=0.15P PS=1.012U PD=2.596U
.ENDS inverter__inv

*** SUBCIRCUIT Repeater__Repeater FROM CELL Repeater:Repeater{lay}
.SUBCKT Repeater__Repeater gnd in out vdd
Xinv@1 gnd in net@7 vdd inverter__inv
Xinv@2 gnd net@7 out vdd inverter__inv
.ENDS Repeater__Repeater

*** TOP LEVEL CELL: Repeater:Repeater_sim{lay}
XRepeater@0 gnd in out vdd Repeater__Repeater

* Spice Code nodes in cell cell 'Repeater:Repeater_sim{lay}'
vdd vdd 0 DC 0.95
vin in 0 DC pwl 10n 0 20n 0.95 50n 0.95 60n 0
cload out 0 250fF
.measure tran tf trig v(out) val=4.5 fall=1 td=8ns targ v(out) val=0.5 fall=1
.measure tran tr trig v(out) val=0.5 rise=1 td=50ns targ v(out) val=4.5 rise=1
.tran 0 100ns
.include C:\Electric\22nm.txt
.END
