*** SPICE deck for cell inv_90nm{sch} from library inverter
*** Created on Thu Jan 02, 2025 17:48:16
*** Last revised on Thu Jan 02, 2025 22:12:49
*** Written on Thu Jan 02, 2025 22:12:53 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: inverter:inv_90nm{sch}
Mnmos@0 out in gnd gnd N L=0.044U W=0.22U
Mpmos@0 vdd in out vdd P L=0.044U W=0.44U

* Spice Code nodes in cell cell 'inverter:inv_90nm{sch}'
vdd vdd 0 DC 0.95
vin in 0 DC pwl 10n 0 20n 0.95 50n 0.95 60n 0
cload out 0 250fF
.measure tran tf trig v(out) val=4.5 fall=1 td=8ns targ v(out) val=0.5 fall=1
.measure tran tr trig v(out) val=0.5 rise=1 td=50ns targ v(out) val=4.5 rise=1
.tran 0 100ns
.include C:\Electric\22nm.txt
.END
