*** SPICE deck for cell 2bit_FA_leftSide_sim{lay} from library 2bit_FA
*** Created on Mon Jan 13, 2025 22:23:11
*** Last revised on Mon Jan 13, 2025 22:34:26
*** Written on Mon Jan 13, 2025 22:34:41 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT _2bit_FA__2bit_FA_leftSide FROM CELL 2bit_FA:2bit_FA_leftSide{lay}
.SUBCKT _2bit_FA__2bit_FA_leftSide A2 A3 B2 B3 c1 c2 G2 G3 gnd P2 P3 s2 s3 vdd
Mnmos@0 gnd b2 net@3 gnd N L=0.044U W=0.22U AS=0.015P AD=0.161P PS=0.352U PD=1.875U
Mnmos@1 net@3 a2 G2 gnd N L=0.044U W=0.22U AS=0.045P AD=0.015P PS=0.689U PD=0.352U
Mnmos@2 net@14 a2 P2 gnd N L=0.044U W=0.44U AS=0.067P AD=0.047P PS=0.858U PD=0.875U
Mnmos@3 P2 net@22 net@14 gnd N L=0.044U W=0.44U AS=0.047P AD=0.067P PS=0.875U PD=0.858U
Mnmos@4 net@14 net@15 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.047P PS=1.875U PD=0.875U
Mnmos@5 gnd b2 net@14 gnd N L=0.044U W=0.44U AS=0.047P AD=0.161P PS=0.875U PD=1.875U
Mnmos@6 gnd a2 net@15 gnd N L=0.044U W=0.44U AS=0.087P AD=0.161P PS=1.584U PD=1.875U
Mnmos@7 net@22 b2 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.087P PS=1.875U PD=1.584U
Mnmos@8 net@64 P2 s2 gnd N L=0.044U W=0.44U AS=0.067P AD=0.047P PS=0.858U PD=0.875U
Mnmos@9 s2 net@71 net@64 gnd N L=0.044U W=0.44U AS=0.047P AD=0.067P PS=0.875U PD=0.858U
Mnmos@10 net@64 net@65 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.047P PS=1.875U PD=0.875U
Mnmos@11 gnd c1 net@64 gnd N L=0.044U W=0.44U AS=0.047P AD=0.161P PS=0.875U PD=1.875U
Mnmos@12 gnd P2 net@65 gnd N L=0.044U W=0.44U AS=0.087P AD=0.161P PS=1.584U PD=1.875U
Mnmos@13 net@71 c1 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.087P PS=1.875U PD=1.584U
Mnmos@14 gnd b3 net@307 gnd N L=0.044U W=0.22U AS=0.015P AD=0.161P PS=0.352U PD=1.875U
Mnmos@15 net@307 a3 G3 gnd N L=0.044U W=0.22U AS=0.045P AD=0.015P PS=0.689U PD=0.352U
Mnmos@16 net@238 a3 P3 gnd N L=0.044U W=0.44U AS=0.067P AD=0.047P PS=0.858U PD=0.875U
Mnmos@17 P3 net@254 net@238 gnd N L=0.044U W=0.44U AS=0.047P AD=0.067P PS=0.875U PD=0.858U
Mnmos@18 net@238 net@249 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.047P PS=1.875U PD=0.875U
Mnmos@19 gnd b3 net@238 gnd N L=0.044U W=0.44U AS=0.047P AD=0.161P PS=0.875U PD=1.875U
Mnmos@20 gnd a3 net@249 gnd N L=0.044U W=0.44U AS=0.087P AD=0.161P PS=1.584U PD=1.875U
Mnmos@21 net@254 b3 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.087P PS=1.875U PD=1.584U
Mnmos@22 net@197 P3 s3 gnd N L=0.044U W=0.44U AS=0.067P AD=0.047P PS=0.858U PD=0.875U
Mnmos@23 s3 net@253 net@197 gnd N L=0.044U W=0.44U AS=0.047P AD=0.067P PS=0.875U PD=0.858U
Mnmos@24 net@197 net@196 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.047P PS=1.875U PD=0.875U
Mnmos@25 gnd c2 net@197 gnd N L=0.044U W=0.44U AS=0.047P AD=0.161P PS=0.875U PD=1.875U
Mnmos@26 gnd P3 net@196 gnd N L=0.044U W=0.44U AS=0.087P AD=0.161P PS=1.584U PD=1.875U
Mnmos@27 net@253 c2 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.087P PS=1.875U PD=1.584U
Mpmos@0 vdd b2 G2 vdd P L=0.044U W=0.44U AS=0.045P AD=0.213P PS=0.689U PD=2.695U
Mpmos@1 G2 a2 vdd vdd P L=0.044U W=0.44U AS=0.213P AD=0.045P PS=2.695U PD=0.689U
Mpmos@2 vdd a2 net@48 vdd P L=0.044U W=0.88U AS=0.053P AD=0.213P PS=1.001U PD=2.695U
Mpmos@3 net@48 net@22 P2 vdd P L=0.044U W=0.88U AS=0.067P AD=0.053P PS=0.858U PD=1.001U
Mpmos@4 P2 net@15 net@51 vdd P L=0.044U W=0.88U AS=0.053P AD=0.067P PS=1.001U PD=0.858U
Mpmos@5 net@51 b2 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.053P PS=2.695U PD=1.001U
Mpmos@6 vdd a2 net@15 vdd P L=0.044U W=0.88U AS=0.087P AD=0.213P PS=1.584U PD=2.695U
Mpmos@7 net@22 b2 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.087P PS=2.695U PD=1.584U
Mpmos@8 vdd P2 net@97 vdd P L=0.044U W=0.88U AS=0.053P AD=0.213P PS=1.001U PD=2.695U
Mpmos@9 net@97 net@71 s2 vdd P L=0.044U W=0.88U AS=0.067P AD=0.053P PS=0.858U PD=1.001U
Mpmos@10 s2 net@65 net@100 vdd P L=0.044U W=0.88U AS=0.053P AD=0.067P PS=1.001U PD=0.858U
Mpmos@11 net@100 c1 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.053P PS=2.695U PD=1.001U
Mpmos@12 vdd P2 net@65 vdd P L=0.044U W=0.88U AS=0.087P AD=0.213P PS=1.584U PD=2.695U
Mpmos@13 net@71 c1 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.087P PS=2.695U PD=1.584U
Mpmos@14 vdd b3 G3 vdd P L=0.044U W=0.44U AS=0.045P AD=0.213P PS=0.689U PD=2.695U
Mpmos@15 G3 a3 vdd vdd P L=0.044U W=0.44U AS=0.213P AD=0.045P PS=2.695U PD=0.689U
Mpmos@16 vdd a3 net@327 vdd P L=0.044U W=0.88U AS=0.053P AD=0.213P PS=1.001U PD=2.695U
Mpmos@17 net@327 net@254 P3 vdd P L=0.044U W=0.88U AS=0.067P AD=0.053P PS=0.858U PD=1.001U
Mpmos@18 P3 net@249 net@331 vdd P L=0.044U W=0.88U AS=0.053P AD=0.067P PS=1.001U PD=0.858U
Mpmos@19 net@331 b3 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.053P PS=2.695U PD=1.001U
Mpmos@20 vdd a3 net@249 vdd P L=0.044U W=0.88U AS=0.087P AD=0.213P PS=1.584U PD=2.695U
Mpmos@21 net@254 b3 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.087P PS=2.695U PD=1.584U
Mpmos@22 vdd P3 net@381 vdd P L=0.044U W=0.88U AS=0.053P AD=0.213P PS=1.001U PD=2.695U
Mpmos@23 net@381 net@253 s3 vdd P L=0.044U W=0.88U AS=0.067P AD=0.053P PS=0.858U PD=1.001U
Mpmos@24 s3 net@196 net@195 vdd P L=0.044U W=0.88U AS=0.053P AD=0.067P PS=1.001U PD=0.858U
Mpmos@25 net@195 c2 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.053P PS=2.695U PD=1.001U
Mpmos@26 vdd P3 net@196 vdd P L=0.044U W=0.88U AS=0.087P AD=0.213P PS=1.584U PD=2.695U
Mpmos@27 net@253 c2 vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.087P PS=2.695U PD=1.584U
.ENDS _2bit_FA__2bit_FA_leftSide

*** TOP LEVEL CELL: 2bit_FA:2bit_FA_leftSide_sim{lay}
X_2bit_FA_@0 A2 A3 B2 B3 c1 c2 G2 G3 gnd P2 P3 s2 s3 vdd _2bit_FA__2bit_FA_leftSide

* Spice Code nodes in cell cell '2bit_FA:2bit_FA_leftSide_sim{lay}'
vdd vdd 0 DC 0.95
* 2-bit input A
va2 A2 0 PWL(0n 0 10n 0 12n 0.95 51n 0.95 53n 0 95n 0 97n 0.95 140n 0.95 142n 0 183n 0 185n 0.95)
va3 A3 0 PWL(0n 0.95 10n 0.95 12n 0 51n 0 53n 0.95 95n 0.95 97n 0 140n 0 142n 0.95 183n 0.95 185n 0)
* 2-bit input B
vb2 B2 0 PWL(0n 0 95n 0 97n 0.95)
vb3 B3 0 PWL(0n 0.95 95n 0.95 97n 0)
vc1 c1 0 DC 0
vc2 c2 0 DC 0
* Transient analysis
.tran 0 200n
* Include model file
.include C:\Electric\22nm.txt
.END
