*** SPICE deck for cell 4bit_FA_block{lay} from library FA_for_CLA
*** Created on Tue Jan 07, 2025 17:49:34
*** Last revised on Fri Jan 10, 2025 21:22:35
*** Written on Fri Jan 10, 2025 21:22:40 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT XOR__XOR FROM CELL XOR:XOR{lay}
.SUBCKT XOR__XOR A B gnd out vdd
Mnmos@0 net@3 A out gnd N L=0.044U W=0.44U AS=0.067P AD=0.047P PS=0.858U PD=0.875U
Mnmos@1 out net@256 net@3 gnd N L=0.044U W=0.44U AS=0.047P AD=0.067P PS=0.875U PD=0.858U
Mnmos@4 net@3 net@199 gnd gnd N L=0.044U W=0.44U AS=0.165P AD=0.047P PS=2.04U PD=0.875U
Mnmos@5 gnd B net@3 gnd N L=0.044U W=0.44U AS=0.047P AD=0.165P PS=0.875U PD=2.04U
Mnmos@7 gnd A net@199 gnd N L=0.044U W=0.44U AS=0.087P AD=0.165P PS=1.584U PD=2.04U
Mnmos@9 net@256 B gnd gnd N L=0.044U W=0.44U AS=0.165P AD=0.087P PS=2.04U PD=1.584U
Mpmos@0 vdd A net@477 vdd P L=0.044U W=0.88U AS=0.053P AD=0.238P PS=1.001U PD=3.196U
Mpmos@1 net@477 net@256 out vdd P L=0.044U W=0.88U AS=0.067P AD=0.053P PS=0.858U PD=1.001U
Mpmos@4 out net@199 net@497 vdd P L=0.044U W=0.88U AS=0.053P AD=0.067P PS=1.001U PD=0.858U
Mpmos@5 net@497 B vdd vdd P L=0.044U W=0.88U AS=0.238P AD=0.053P PS=3.196U PD=1.001U
Mpmos@6 vdd A net@199 vdd P L=0.044U W=0.88U AS=0.087P AD=0.238P PS=1.584U PD=3.196U
Mpmos@7 net@256 B vdd vdd P L=0.044U W=0.88U AS=0.238P AD=0.087P PS=3.196U PD=1.584U
.ENDS XOR__XOR

*** SUBCIRCUIT NAND__nand FROM CELL NAND:nand{lay}
.SUBCKT NAND__nand A B gnd out vdd
Mnmos@0 gnd B net@45 gnd N L=0.044U W=0.22U AS=0.015P AD=0.106P PS=0.352U PD=2.288U
Mnmos@1 net@45 A out gnd N L=0.044U W=0.22U AS=0.047P AD=0.015P PS=0.704U PD=0.352U
Mpmos@0 vdd B out vdd P L=0.044U W=0.44U AS=0.047P AD=0.106P PS=0.704U PD=1.969U
Mpmos@1 out A vdd vdd P L=0.044U W=0.44U AS=0.106P AD=0.047P PS=1.969U PD=0.704U
.ENDS NAND__nand

*** SUBCIRCUIT FA_for_CLA__FA FROM CELL FA_for_CLA:FA{lay}
.SUBCKT FA_for_CLA__FA A B Cin G gnd P Sum vdd
XXOR@0 a b gnd P vdd XOR__XOR
XXOR@1 P cin gnd Sum vdd XOR__XOR
Xnand@0 a b gnd G vdd NAND__nand
.ENDS FA_for_CLA__FA

*** SUBCIRCUIT FA_for_CLA__4bit_FA FROM CELL FA_for_CLA:4bit_FA{lay}
.SUBCKT FA_for_CLA__4bit_FA A0 A1 A2 A3 B0 B1 B2 B3 c-1 c0 c1 c2 G0 G1 G2 G3 gnd P0 P1 P2 P3 s0 s1 s2 s3 vdd
XFA@0 A0 B0 c-1 G0 gnd P0 s0 vdd FA_for_CLA__FA
XFA@1 A1 B1 c0 G1 gnd P1 s1 vdd FA_for_CLA__FA
XFA@2 A2 B2 c1 G2 gnd P2 s2 vdd FA_for_CLA__FA
XFA@3 A3 B3 c2 G3 gnd P3 s3 vdd FA_for_CLA__FA
.ENDS FA_for_CLA__4bit_FA

*** TOP LEVEL CELL: FA_for_CLA:4bit_FA_block{lay}
X_4bit_FA@0 A0 A1 A2 A3 B0 B1 B2 B3 c-1 c0 c1 c2 G0 G1 G2 G3 gnd P0 P1 P2 P3 s0 s1 s2 s3 vdd FA_for_CLA__4bit_FA

* Spice Code nodes in cell cell 'FA_for_CLA:4bit_FA_block{lay}'
* 4-bit Carry Look-Ahead Adder Simulation
* Power supply
vdd vdd 0 DC 0.95
cload0 s0 0 50fF
cload1 s1 0 50fF
cload2 s2 0 50fF
cload3 s3 0 50fF
* 4-bit input A
va0 A0 0 PWL(0n 0 10n 0 12n 0.95 51n 0.95 53n 0 95n 0 97n 0.95 140n 0.95 142n 0 183n 0 185n 0.95)
va1 A1 0 PWL(0n 0.95 10n 0.95 12n 0 51n 0 53n 0.95 95n 0.95 97n 0 140n 0 142n 0.95 183n 0.95 185n 0)
va2 A2 0 PWL(0n 0 10n 0 12n 0.95 51n 0.95 53n 0 95n 0 97n 0.95 140n 0.95 142n 0 183n 0 185n 0.95)
va3 A3 0 PWL(0n 0.95 10n 0.95 12n 0 51n 0 53n 0.95 95n 0.95 97n 0 140n 0 142n 0.95 183n 0.95 185n 0)
* 4-bit input B
vb0 B0 0 PWL(0n 0 95n 0 97n 0.95)
vb1 B1 0 PWL(0n 0.95 95n 0.95 97n 0)
vb2 B2 0 PWL(0n 0 95n 0 97n 0.95)
vb3 B3 0 PWL(0n 0.95 95n 0.95 97n 0)
* Initial carry-in C0
vc-1 c-1 0 DC 0.95
vc0 c0 0 DC 0
vc1 c1 0 DC 0
vc2 c2 0 DC 0.95
* Clock signal
vclk clk 0 PWL(0n 0 20n 0 22n 0.95 42n 0.95 44n 0 64n 0 66n 0.95 86n 0.95 88n 0 108n 0 110n 0.95 130n 0.95 132n 0 152n 0 154n 0.95 174n 0.95 176n 0 196n 0 198n 0.95)
* Transient analysis
.tran 0 200n
* Include model file
.include C:\Electric\22nm.txt
.END
