*** SPICE deck for cell nand{lay} from library NAND
*** Created on Sat Nov 09, 2024 20:34:09
*** Last revised on Thu Jan 02, 2025 14:40:47
*** Written on Thu Jan 02, 2025 14:40:53 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: NAND:nand{lay}
Mnmos@0 gnd B net@45 gnd N L=0.6U W=3U AS=2.7P AD=19.8P PS=4.8U PD=31.2U
Mnmos@1 net@45 A out gnd N L=0.6U W=3U AS=8.7P AD=2.7P PS=9.6U PD=4.8U
Mpmos@0 vdd B out vdd P L=0.6U W=6U AS=8.7P AD=19.8P PS=9.6U PD=26.85U
Mpmos@1 out A vdd vdd P L=0.6U W=6U AS=19.8P AD=8.7P PS=26.85U PD=9.6U

* Spice Code nodes in cell cell 'NAND:nand{lay}'
vdd vdd 0 DC 5
va A 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb B 0 DC pwl 10n 0 20n 5 100n 5 110n 0
.measure tran tf trig v(out) val=4.5 fall=1 td=4ns trag v(out) val=0.5 fall=1
.measure tran tr trig v(out) val=0.5 rise=1 td=4ns trag v(out) val=4.5 rise=1
.tran 200n
.include C:\Electric\C5_models.txt
.END
