*** SPICE deck for cell XOR_sim{lay} from library XOR
*** Created on Sun Nov 10, 2024 12:25:45
*** Last revised on Thu Jan 02, 2025 14:34:45
*** Written on Thu Jan 02, 2025 14:34:51 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT XOR__XOR FROM CELL XOR:XOR{lay}
.SUBCKT XOR__XOR A B gnd out vdd
Mnmos@0 net@3 A out gnd N L=0.6U W=3U AS=6.638P AD=4.725P PS=7.275U PD=7.65U
Mnmos@1 out net@202 net@3 gnd N L=0.6U W=3U AS=4.725P AD=6.638P PS=7.65U PD=7.275U
Mnmos@4 net@3 net@191 gnd gnd N L=0.6U W=3U AS=25.988P AD=4.725P PS=23.325U PD=7.65U
Mnmos@5 gnd B net@3 gnd N L=0.6U W=3U AS=4.725P AD=25.988P PS=7.65U PD=23.325U
Mnmos@7 gnd A net@191 gnd N L=0.6U W=3U AS=8.325P AD=25.988P PS=12.75U PD=23.325U
Mnmos@9 net@202 B gnd gnd N L=0.6U W=3U AS=25.988P AD=8.1P PS=23.325U PD=12.6U
Mpmos@0 vdd A net@236 vdd P L=0.6U W=6U AS=4.5P AD=33.75P PS=7.5U PD=31.875U
Mpmos@1 net@236 net@202 out vdd P L=0.6U W=6U AS=6.638P AD=4.5P PS=7.275U PD=7.5U
Mpmos@4 out net@191 net@240 vdd P L=0.6U W=6U AS=5.4P AD=6.638P PS=7.8U PD=7.275U
Mpmos@5 net@240 B vdd vdd P L=0.6U W=6U AS=33.75P AD=5.4P PS=31.875U PD=7.8U
Mpmos@6 vdd A net@191 vdd P L=0.6U W=6U AS=8.325P AD=33.75P PS=12.75U PD=31.875U
Mpmos@7 net@202 B vdd vdd P L=0.6U W=6U AS=33.75P AD=8.1P PS=31.875U PD=12.6U
.ENDS XOR__XOR

*** TOP LEVEL CELL: XOR:XOR_sim{lay}
XXOR@0 A B gnd out vdd XOR__XOR

* Spice Code nodes in cell cell 'XOR:XOR_sim{lay}'
vdd vdd 0 DC 5
va A 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb B 0 DC pwl 10n 0 20n 5 100n 5 110n 0
.tran 200n
.include C:\Electric\C5_models.txt
.END
