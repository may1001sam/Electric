*** SPICE deck for cell FA_new_sim{lay} from library FA_new
*** Created on Mon Jan 13, 2025 18:06:10
*** Last revised on Mon Jan 13, 2025 21:01:26
*** Written on Mon Jan 13, 2025 21:01:37 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT FA_new__FA_new FROM CELL FA_new:FA_new{lay}
.SUBCKT FA_new__FA_new A B Cin G gnd P Sum vdd
Mnmos@12 gnd b net@157 gnd N L=0.044U W=0.22U AS=0.015P AD=0.161P PS=0.352U PD=1.875U
Mnmos@13 net@157 a G gnd N L=0.044U W=0.22U AS=0.045P AD=0.015P PS=0.689U PD=0.352U
Mnmos@14 net@175 a P gnd N L=0.044U W=0.44U AS=0.067P AD=0.047P PS=0.858U PD=0.875U
Mnmos@15 P net@183 net@175 gnd N L=0.044U W=0.44U AS=0.047P AD=0.067P PS=0.875U PD=0.858U
Mnmos@16 net@175 net@176 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.047P PS=1.875U PD=0.875U
Mnmos@17 gnd b net@175 gnd N L=0.044U W=0.44U AS=0.047P AD=0.161P PS=0.875U PD=1.875U
Mnmos@18 gnd a net@176 gnd N L=0.044U W=0.44U AS=0.087P AD=0.161P PS=1.584U PD=1.875U
Mnmos@19 net@183 b gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.087P PS=1.875U PD=1.584U
Mnmos@20 net@251 P Sum gnd N L=0.044U W=0.44U AS=0.067P AD=0.047P PS=0.858U PD=0.875U
Mnmos@21 Sum net@259 net@251 gnd N L=0.044U W=0.44U AS=0.047P AD=0.067P PS=0.875U PD=0.858U
Mnmos@22 net@251 net@252 gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.047P PS=1.875U PD=0.875U
Mnmos@23 gnd cin net@251 gnd N L=0.044U W=0.44U AS=0.047P AD=0.161P PS=0.875U PD=1.875U
Mnmos@24 gnd P net@252 gnd N L=0.044U W=0.44U AS=0.087P AD=0.161P PS=1.584U PD=1.875U
Mnmos@25 net@259 cin gnd gnd N L=0.044U W=0.44U AS=0.161P AD=0.087P PS=1.875U PD=1.584U
Mpmos@12 vdd b G vdd P L=0.044U W=0.44U AS=0.045P AD=0.213P PS=0.689U PD=2.695U
Mpmos@13 G a vdd vdd P L=0.044U W=0.44U AS=0.213P AD=0.045P PS=2.695U PD=0.689U
Mpmos@14 vdd a net@216 vdd P L=0.044U W=0.88U AS=0.053P AD=0.213P PS=1.001U PD=2.695U
Mpmos@15 net@216 net@183 P vdd P L=0.044U W=0.88U AS=0.067P AD=0.053P PS=0.858U PD=1.001U
Mpmos@16 P net@176 net@219 vdd P L=0.044U W=0.88U AS=0.053P AD=0.067P PS=1.001U PD=0.858U
Mpmos@17 net@219 b vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.053P PS=2.695U PD=1.001U
Mpmos@18 vdd a net@176 vdd P L=0.044U W=0.88U AS=0.087P AD=0.213P PS=1.584U PD=2.695U
Mpmos@19 net@183 b vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.087P PS=2.695U PD=1.584U
Mpmos@20 vdd P net@292 vdd P L=0.044U W=0.88U AS=0.053P AD=0.213P PS=1.001U PD=2.695U
Mpmos@21 net@292 net@259 Sum vdd P L=0.044U W=0.88U AS=0.067P AD=0.053P PS=0.858U PD=1.001U
Mpmos@22 Sum net@252 net@295 vdd P L=0.044U W=0.88U AS=0.053P AD=0.067P PS=1.001U PD=0.858U
Mpmos@23 net@295 cin vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.053P PS=2.695U PD=1.001U
Mpmos@24 vdd P net@252 vdd P L=0.044U W=0.88U AS=0.087P AD=0.213P PS=1.584U PD=2.695U
Mpmos@25 net@259 cin vdd vdd P L=0.044U W=0.88U AS=0.213P AD=0.087P PS=2.695U PD=1.584U
.ENDS FA_new__FA_new

*** TOP LEVEL CELL: FA_new:FA_new_sim{lay}
XFA_new@2 A B Cin G gnd P Sum vdd FA_new__FA_new

* Spice Code nodes in cell cell 'FA_new:FA_new_sim{lay}'
* 4-bit Carry Look-Ahead Adder Simulation
* Power supply
vdd vdd 0 DC 0.95
va A 0 PWL(0n 0 10n 0 12n 0.95 51n 0.95 53n 0 95n 0 97n 0.95 140n 0.95 142n 0 183n 0 185n 0.95)
vb B 0 PWL(0n 0 95n 0 97n 0.95)
vcin Cin 0 DC 0.95
* Transient analysis
.tran 0 200n
* Include model file
.include C:\Electric\22nm.txt
.END
