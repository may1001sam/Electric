*** SPICE deck for cell nand{sch} from library NAND
*** Created on Sat Nov 09, 2024 14:22:29
*** Last revised on Thu Jan 02, 2025 22:43:31
*** Written on Thu Jan 02, 2025 22:43:34 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: NAND:nand{sch}
Mnmos@0 out A net@11 gnd N L=0.044U W=0.22U
Mnmos@1 net@11 B gnd gnd N L=0.044U W=0.33U
Mpmos@1 vdd A out vdd P L=0.044U W=0.44U
Mpmos@2 vdd B out vdd P L=0.044U W=0.44U

* Spice Code nodes in cell cell 'NAND:nand{sch}'
vdd vdd 0 DC 0.95
va A 0 DC pwl 10n 0 20n 0.95 50n 0.95 60n 0 90n 0 100n 0.95 130n 0.95 140n 0 170n 0 180n 0.95
vb B 0 DC pwl 10n 0 20n 0.95 100n 0.95 110n 0
.tran 200n
.include C:\Electric\22nm.txt
.END
